module and_gate (
    input logic a, b,
    output logic y
);
    assign y = a && b; // Using logical AND operator
endmodule

